//AND logic
module AND_logic(
    input branch,zero,
    output and_out
    );
    assign and_out = branch & zero;
endmodule
